module add ;
